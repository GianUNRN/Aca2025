module button (
    input logic bt,
    output logic out_bt
);
    assign out_bt = bt;
endmodule