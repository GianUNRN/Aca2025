module switches (
    input logic [7:0] sw,
    output logic [7:0] decoded_swithces
);
    assign decoded_swithces = sw;
endmodule